library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.numeric_std.all;

package registers is
	type reg_array is array(31 downto 0) of std_logic_vector (31 downto 0); 
end package registers;
package body registers is
end package body registers;